module display #(parameter NUM_SEGMENTS, parameter ASCII_LEN) (ascii, HEX);
    input  logic [   ASCII_LEN-1:0] ascii;
    output logic [NUM_SEGMENTS-1:0] HEX;

    always_comb begin
        HEX = 8'b11111111;  // space
        case (ascii)
            8'h20  : HEX = 8'b11111111;  // space
            8'h21  : HEX = 8'b01111001;  // !
            8'h22  : HEX = 8'b11011101;  // "
            8'h23  : HEX = 8'b10000001;  // #
            8'h24  : HEX = 8'b10010010;  // $
            8'h25  : HEX = 8'b00101101;  // %
            8'h26  : HEX = 8'b10111001;  // &
            8'h27  : HEX = 8'b11011111;  // '
            8'h28  : HEX = 8'b11010110;  // (
            8'h29  : HEX = 8'b11110100;  // )
            8'h2a  : HEX = 8'b11011110;  // *
            8'h2b  : HEX = 8'b10001111;  // +
            8'h2c  : HEX = 8'b11101111;  // ,
            8'h2d  : HEX = 8'b10111111;  // -
            8'h2e  : HEX = 8'b01111111;  // .
            8'h2f  : HEX = 8'b10101101;  // /
            8'h30  : HEX = 8'b11000000;  // 0
            8'h31  : HEX = 8'b11111001;  // 1
            8'h32  : HEX = 8'b10100100;  // 2
            8'h33  : HEX = 8'b10110000;  // 3
            8'h34  : HEX = 8'b10011001;  // 4
            8'h35  : HEX = 8'b10010010;  // 5
            8'h36  : HEX = 8'b10000010;  // 6
            8'h37  : HEX = 8'b11111000;  // 7
            8'h38  : HEX = 8'b10000000;  // 8
            8'h39  : HEX = 8'b10010000;  // 9
            8'h3a  : HEX = 8'b11110110;  // :
            8'h3b  : HEX = 8'b11110010;  // ;
            8'h3c  : HEX = 8'b10011110;  // <
            8'h3d  : HEX = 8'b10110111;  // =
            8'h3e  : HEX = 8'b10111100;  // >
            8'h3f  : HEX = 8'b00101100;  // ?
            8'h40  : HEX = 8'b10100000;  // @
            8'h41  : HEX = 8'b10001000;  // A
            8'h42  : HEX = 8'b10000011;  // B
            8'h43  : HEX = 8'b11000110;  // C
            8'h44  : HEX = 8'b10100001;  // D
            8'h45  : HEX = 8'b10000110;  // E
            8'h46  : HEX = 8'b10001110;  // F
            8'h47  : HEX = 8'b11000010;  // G
            8'h48  : HEX = 8'b10001001;  // H
            8'h49  : HEX = 8'b11001111;  // I
            8'h4a  : HEX = 8'b11100001;  // J
            8'h4b  : HEX = 8'b10001010;  // K
            8'h4c  : HEX = 8'b11000111;  // L
            8'h4d  : HEX = 8'b11101010;  // M
            8'h4e  : HEX = 8'b11001000;  // N
            8'h4f  : HEX = 8'b11000000;  // O
            8'h50  : HEX = 8'b10001100;  // P
            8'h51  : HEX = 8'b10010100;  // Q
            8'h52  : HEX = 8'b11001100;  // R
            8'h53  : HEX = 8'b10010010;  // S
            8'h54  : HEX = 8'b10000111;  // T
            8'h55  : HEX = 8'b11000001;  // U
            8'h56  : HEX = 8'b11000001;  // V
            8'h57  : HEX = 8'b11010101;  // W
            8'h58  : HEX = 8'b10001001;  // X
            8'h59  : HEX = 8'b10010001;  // Y
            8'h5a  : HEX = 8'b10100100;  // Z
            8'h5b  : HEX = 8'b11000110;  // [
            8'h5c  : HEX = 8'b10011011;  // \
            8'h5d  : HEX = 8'b11110000;  // ]
            8'h5e  : HEX = 8'b11011100;  // ^
            8'h5f  : HEX = 8'b11110111;  // _
            8'h60  : HEX = 8'b11111101;  // `
            8'h61  : HEX = 8'b10100000;  // a
            8'h62  : HEX = 8'b10000011;  // b
            8'h63  : HEX = 8'b10100111;  // c
            8'h64  : HEX = 8'b10100001;  // d
            8'h65  : HEX = 8'b10000100;  // e
            8'h66  : HEX = 8'b10001110;  // f
            8'h67  : HEX = 8'b10010000;  // g
            8'h68  : HEX = 8'b10001011;  // h
            8'h69  : HEX = 8'b11101111;  // i
            8'h6a  : HEX = 8'b11110011;  // j
            8'h6b  : HEX = 8'b10001010;  // k
            8'h6c  : HEX = 8'b11001111;  // l
            8'h6d  : HEX = 8'b11101011;  // m
            8'h6e  : HEX = 8'b10101011;  // n
            8'h6f  : HEX = 8'b10100011;  // o
            8'h70  : HEX = 8'b10001100;  // p
            8'h71  : HEX = 8'b10011000;  // q
            8'h72  : HEX = 8'b10101111;  // r
            8'h73  : HEX = 8'b10010010;  // s
            8'h74  : HEX = 8'b10000111;  // t
            8'h75  : HEX = 8'b11100011;  // u
            8'h76  : HEX = 8'b11100011;  // v
            8'h77  : HEX = 8'b11101011;  // /
            8'h78  : HEX = 8'b10001001;  // x
            8'h79  : HEX = 8'b10010001;  // y
            8'h7a  : HEX = 8'b10100100;  // z
            8'h7b  : HEX = 8'b10111001;  // {
            8'h7c  : HEX = 8'b11001111;  // |
            8'h7d  : HEX = 8'b10001111;  // }
            8'h7e  : HEX = 8'b11111110;  // ~
            default: ;
        endcase
    end
endmodule
